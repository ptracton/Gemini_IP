/*
 * File: gpio_agent.sv
 * Description: GPIO Agent
 */

class gpio_agent extends uvm_agent;
    `uvm_component_utils(gpio_agent)

    gpio_driver    driver;
    uvm_sequencer #(gpio_seq_item) sequencer;
    gpio_monitor   monitor;

    function new(string name, uvm_component parent);
        super.new(name, parent);
    endfunction

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        monitor = gpio_monitor::type_id::create("monitor", this);
        if (get_is_active() == UVM_ACTIVE) begin
            driver = gpio_driver::type_id::create("driver", this);
            sequencer = uvm_sequencer#(gpio_seq_item)::type_id::create("sequencer", this);
        end
    endfunction

    function void connect_phase(uvm_phase phase);
        if (get_is_active() == UVM_ACTIVE) begin
            driver.seq_item_port.connect(sequencer.seq_item_export);
        end
    endfunction

endclass
