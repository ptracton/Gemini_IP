
// Interfaces and Packages
`include "apb_if.sv"
`include "axi_if.sv"
`include "wb_if.sv"
`include "agents/uart_agent/uart_if.sv"

`include "apb_agent_pkg.sv"
`include "axi_agent_pkg.sv"
`include "wb_agent_pkg.sv"
`include "agents/uart_agent/uart_agent_pkg.sv"
`include "env/uart_env_pkg.sv"
`include "tests/uart_test_pkg.sv"

// DUT files and TB files are compiled separately
