/*
 * File: gpio_agent_pkg.sv
 * Description: GPIO Agent Package
 */

package gpio_agent_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "gpio_seq_item.sv"
    `include "gpio_driver.sv"
    `include "gpio_monitor.sv"
    `include "gpio_agent.sv"

endpackage
