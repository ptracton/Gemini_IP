/*
 * File: bus_matrix_agent_pkg.sv
 * Description: UVM Package for Timer specific IO Agent
 */
package bus_matrix_agent_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "bus_matrix_seq_item.sv"
    `include "bus_matrix_driver.sv"
    `include "bus_matrix_monitor.sv"
    `include "bus_matrix_agent.sv"

endpackage
