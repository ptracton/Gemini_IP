/*
 * File: ahb_agent_pkg.sv
 * Description: AHB Agent Package
 */

package ahb_agent_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "ahb_seq_item.sv"
    `include "ahb_seq.sv"
    `include "ahb_driver.sv"
    `include "ahb_slave_driver.sv"
    `include "ahb_monitor.sv"
    `include "ahb_agent.sv"

endpackage
