`ifndef SPI_AGENT_SV
`define SPI_AGENT_SV

`include "spi_seq_item.sv"
`include "spi_driver.sv"
`include "spi_monitor.sv"
`include "spi_sequencer.sv"

class spi_agent extends uvm_agent;
  `uvm_component_utils(spi_agent)

  spi_driver    driver;
  spi_monitor   monitor;
  spi_sequencer sequencer;

  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    monitor = spi_monitor::type_id::create("monitor", this);
    if (get_is_active() == UVM_ACTIVE) begin
      driver = spi_driver::type_id::create("driver", this);
      sequencer = spi_sequencer::type_id::create("sequencer", this);
    end
  endfunction

  function void connect_phase(uvm_phase phase);
    if (get_is_active() == UVM_ACTIVE) begin
      driver.seq_item_port.connect(sequencer.seq_item_export);
    end
  endfunction

endclass

`endif
