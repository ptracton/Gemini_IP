`timescale 1ps / 1ps
module glbl;
  wire GSR = 0;
  wire GTS = 0;
endmodule
