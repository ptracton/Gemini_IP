package bus_matrix_seq_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    import axi_agent_pkg::*;
    import ahb_agent_pkg::*;
    import wb_agent_pkg::*;
    // import bus_matrix_env_pkg::*; // Avoid circular if env imports seq logic? usually env imports agents. 
    
    `include "bus_matrix_sequences.sv"
endpackage
