module bus_matrix_apb_vhdl_binds;
    bind bus_matrix_apb apb_props props_apb (
        .pclk(pclk),
        .presetn(presetn),
        .psel(psel),
        .penable(penable),
        .pwrite(pwrite),
        .paddr(paddr),
        .pwdata(pwdata),
        .pready(pready),
        .prdata(prdata),
        .pslverr(pslverr)
    );
endmodule
