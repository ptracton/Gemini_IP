import bus_matrix_pkg::*;

// -----------------------------------------------------------------------------
// File: bus_matrix_ahb.sv
// Module: bus_matrix_ahb
// Description:
//   AHB-Lite Wrapper for the Bus Matrix.
//   Adapts AHB-Lite protocol (Address Phase, Data Phase, HREADY) to the core
//   matrix logic. Handles HREADYOUT generation and stalling during arbitration.
//
// Parameters:
//   - N_MASTERS, M_SLAVES: Dimensions of the matrix.
//   - DATA_WIDTH, ADDR_WIDTH: Bus widths.
//   - REGION_MAP_FLAT: Memory map configuration.
//   - MASTER_SECURE_MASK: Static security attribute (if HPROT not used/overridden).
//
// Signals:
//   Standard AHB-Lite interfaces (HADDR, HTRANS, HWRITE, HWDATA, HRDATA, etc.)
//   for Master Ports and Slave Ports.
//   Special attention to HREADY (Input) vs HREADYOUT (Output) muxing.
// -----------------------------------------------------------------------------
module bus_matrix_ahb #(
    parameter int N_MASTERS = 2,
    parameter int M_SLAVES = 2,
    parameter int DATA_WIDTH = 32,
    parameter int ADDR_WIDTH = 32,
    parameter logic [M_SLAVES*66-1:0] REGION_MAP_FLAT = '0,
    parameter bit USE_DEFAULT_SLAVE = 0,
    parameter int DEFAULT_SLAVE_INDEX = 0,
    parameter bit INPUT_PIPE_STAGES = 0,
    parameter bit OUTPUT_PIPE_STAGES = 0
)(
    input logic HCLK,
    input logic HRESETn,
    
    // Check bus_matrix_pkg for definitions
    
    // Master Interfaces (Slave Ports on Matrix)
    input  logic [N_MASTERS-1:0]                  HSEL_i,      // From Master (actually generated by interconnect usually, but here inputs)
    // Actually, normally specific masters drive Address, Trans, etc. HSEL is derived.
    // For a matrix, masters drive transfers. The matrix IS the HSEL generator.
    // So Masters allow:
    input  logic [N_MASTERS*ADDR_WIDTH-1:0]       HADDR_i,
    input  logic [N_MASTERS*2-1:0]                HTRANS_i,
    input  logic [N_MASTERS-1:0]                  HWRITE_i,
    input  logic [N_MASTERS*3-1:0]                HSIZE_i,
    input  logic [N_MASTERS*3-1:0]                HBURST_i,
    input  logic [N_MASTERS*4-1:0]                HPROT_i,
    input  logic [N_MASTERS*DATA_WIDTH-1:0]       HWDATA_i,
    // Return path to Masters
    output logic [N_MASTERS-1:0]                  HREADYOUT_o, // To Master
    output logic [N_MASTERS*2-1:0]                HRESP_o,
    output logic [N_MASTERS*DATA_WIDTH-1:0]       HRDATA_o,
    
    // Slave Interfaces (Master Ports on Matrix)
    // To Slaves
    output logic [M_SLAVES-1:0]                   HSEL_o,      // To Slave
    output logic [M_SLAVES*ADDR_WIDTH-1:0]        HADDR_o,
    output logic [M_SLAVES*2-1:0]                 HTRANS_o,
    output logic [M_SLAVES-1:0]                   HWRITE_o,
    output logic [M_SLAVES*3-1:0]                 HSIZE_o,
    output logic [M_SLAVES*3-1:0]                 HBURST_o,
    output logic [M_SLAVES*4-1:0]                 HPROT_o,
    output logic [M_SLAVES*DATA_WIDTH-1:0]        HWDATA_o,
    // From Slaves
    input  logic [M_SLAVES-1:0]                   HREADY_i,    // From Slave
    input  logic [M_SLAVES*2-1:0]                 HRESP_i,
    input  logic [M_SLAVES*DATA_WIDTH-1:0]        HRDATA_i
);

    import bus_matrix_pkg::*;

    // ---------------------------------------------------------
    // 1. Decoder Stage (Address Phase)
    // ---------------------------------------------------------
    logic [N_MASTERS-1:0][M_SLAVES-1:0] master_req_matrix;
    logic [N_MASTERS-1:0]               master_decode_err;
    
    genvar m, s;
    generate
        for (m = 0; m < N_MASTERS; m++) begin : GEN_DECODERS
            logic [ADDR_WIDTH-1:0] m_adr;
            logic [1:0]            m_trans;
            assign m_adr   = HADDR_i[m*ADDR_WIDTH +: ADDR_WIDTH];
            assign m_trans = HTRANS_i[m*2 +: 2];
            
            logic [M_SLAVES-1:0] slave_sel;
            logic internal_err;
            
            bus_matrix_decoder #(
                .M_SLAVES(M_SLAVES),
                .ADDR_WIDTH(ADDR_WIDTH),
                .REGION_MAP_FLAT(REGION_MAP_FLAT),
                .USE_DEFAULT_SLAVE(USE_DEFAULT_SLAVE),
                .DEFAULT_SLAVE_INDEX(DEFAULT_SLAVE_INDEX)
            ) u_dec (
                .addr_i(m_adr),
                .valid_i(m_trans[1]), 
                .secure_i(HPROT_i[m*4 + 1]), // HPROT[1] is 'Non-Secure' usually, so secure = !HPROT[1] ? Or typical 1=Privileged. 
                                             // Standard AHB5: HPROT[1] = Non-Secure. 0=Secure, 1=Non-Secure.
                                             // Decoder expects secure_i=1 for Secure. So secure_i = !HPROT[1].
                .slave_sel_o(slave_sel),
                .dec_error_o(internal_err), // Combined decode error
                .sec_error_o() // We can OR this with dec_error for now or handle distinct HRESP
            );
            
            for (s = 0; s < M_SLAVES; s++) begin
                 assign master_req_matrix[m][s] = slave_sel[s];
            end
            assign master_decode_err[m] = internal_err; // Simplified error handling
        end
    endgenerate

    // ---------------------------------------------------------
    // 2. Arbiter Stage (Address Phase)
    // ---------------------------------------------------------
    logic [M_SLAVES-1:0][N_MASTERS-1:0] slave_req_vector;
    logic [M_SLAVES-1:0][N_MASTERS-1:0] slave_gnt_vector_addr; // Grant for Address Phase
    
    generate
        for (s = 0; s < M_SLAVES; s++) begin
            for (m = 0; m < N_MASTERS; m++) begin
                assign slave_req_vector[s][m] = master_req_matrix[m][s];
            end
        end
    endgenerate

    generate
        for (s = 0; s < M_SLAVES; s++) begin : GEN_ARBITERS
            // Need to hold grant if HREADY is low (stall) or for burst lock (omitted for simplicity here)
            // Just handling HREADY stall: Update grant only when HREADY is high?
            // Actually, arbiter runs combinatorially. We register the result.
            
            bus_matrix_arbiter #(
                .N_REQ(N_MASTERS),
                .SCHEME(0) 
            ) u_arb (
                .clk(HCLK),
                .rst_n(HRESETn),
                .req_i(slave_req_vector[s]),
                .hold_i(!HREADY_i[s]), // Hold arbitration if slave is not ready
                .gnt_o(slave_gnt_vector_addr[s])
            );
        end
    endgenerate
    
    // ---------------------------------------------------------
    // 3. Pipeline Register (Address -> Data Phase Grant)
    // ---------------------------------------------------------
    logic [M_SLAVES-1:0][N_MASTERS-1:0] slave_gnt_vector_data;
    
    always_ff @(posedge HCLK or negedge HRESETn) begin
        if (!HRESETn) begin
            slave_gnt_vector_data <= '0;
        end else begin
            for (int i = 0; i < M_SLAVES; i++) begin
                if (HREADY_i[i]) begin
                     slave_gnt_vector_data[i] <= slave_gnt_vector_addr[i];
                end
            end
        end
    end

    // Transposed Grant Vectors for Master-centric logic
    // [N_MASTERS][M_SLAVES]
    logic [N_MASTERS-1:0][M_SLAVES-1:0] master_gnt_vector_addr;
    logic [N_MASTERS-1:0][M_SLAVES-1:0] master_gnt_vector_data;
    
    generate
        for (m = 0; m < N_MASTERS; m++) begin
            for (s = 0; s < M_SLAVES; s++) begin
                assign master_gnt_vector_addr[m][s] = slave_gnt_vector_addr[s][m];
                assign master_gnt_vector_data[m][s] = slave_gnt_vector_data[s][m];
            end
        end
    endgenerate

    // ---------------------------------------------------------
    // 4. Muxing: Address Phase (Master -> Slave)
    // ---------------------------------------------------------
    generate
        for (s = 0; s < M_SLAVES; s++) begin : GEN_SLAVE_ADDR_MUX
            always_comb begin
                // Defaults
                HSEL_o[s]   = 1'b0;
                HADDR_o[s*ADDR_WIDTH +: ADDR_WIDTH] = '0;
                HTRANS_o[s*2 +: 2] = 2'b00; // IDLE
                HWRITE_o[s] = 1'b0;
                HSIZE_o[s*3 +: 3] = 3'b000;
                HBURST_o[s*3 +: 3] = 3'b000;
                HPROT_o[s*4 +: 4] = 4'b0000;
                
                for (int i = 0; i < N_MASTERS; i++) begin
                    if (slave_gnt_vector_addr[s][i]) begin
                        HSEL_o[s]   = 1'b1; // Select the slave
                        HADDR_o[s*ADDR_WIDTH +: ADDR_WIDTH] = HADDR_i[i*ADDR_WIDTH +: ADDR_WIDTH];
                        HTRANS_o[s*2 +: 2] = HTRANS_i[i*2 +: 2];
                        HWRITE_o[s] = HWRITE_i[i];
                        HSIZE_o[s*3 +: 3] = HSIZE_i[i*3 +: 3];
                        HBURST_o[s*3 +: 3] = HBURST_i[i*3 +: 3];
                        HPROT_o[s*4 +: 4] = HPROT_i[i*4 +: 4];
                    end
                end
            end
        end
    endgenerate

    // ---------------------------------------------------------
    // 5. Muxing: Data Phase (Master -> Slave : HWDATA)
    // ---------------------------------------------------------
    generate
        for (s = 0; s < M_SLAVES; s++) begin : GEN_SLAVE_DATA_MUX
            always_comb begin
                HWDATA_o[s*DATA_WIDTH +: DATA_WIDTH] = '0;
                for (int i = 0; i < N_MASTERS; i++) begin
                    // Data steering based on Data Phase Grant
                    if (slave_gnt_vector_data[s][i]) begin
                        HWDATA_o[s*DATA_WIDTH +: DATA_WIDTH] = HWDATA_i[i*DATA_WIDTH +: DATA_WIDTH];
                    end
                end
            end
        end
    endgenerate

    // ---------------------------------------------------------
    // 6. Return Path Muxing (Slave -> Master : HRDATA, HRESP, HREADY)
    // ---------------------------------------------------------
    generate
        for (m = 0; m < N_MASTERS; m++) begin : GEN_MASTER_MUX
            always_comb begin
                // Defaults
                HRDATA_o[m*DATA_WIDTH +: DATA_WIDTH] = '0;
                HRESP_o[m*2 +: 2] = 2'b00; // OKAY
                HREADYOUT_o[m] = 1'b1;
                
                if (master_decode_err[m]) begin
                     // Error response logic for unmapped address
                     HRESP_o[m*2 +: 2] = 2'b01; // ERROR
                end else begin
                    // Mux based on which slave this master was communicating with in the data phase
                    // Using transposed vector: master_gnt_vector_data[m] is [M_SLAVES-1:0]
                    // We iterate over slaves 'i'.
                    for (int i = 0; i < M_SLAVES; i++) begin
                        if (master_gnt_vector_data[m][i]) begin
                             HRDATA_o[m*DATA_WIDTH +: DATA_WIDTH] = HRDATA_i[i*DATA_WIDTH +: DATA_WIDTH];
                             HRESP_o[m*2 +: 2] = HRESP_i[i*2 +: 2];
                             HREADYOUT_o[m] = HREADY_i[i];
                        end
                    end
                    
                    // Address Phase Stalling (Arbitration Latency)
                    if (HTRANS_i[m*2 + 1]) begin 
                        // Check if any slave granted address phase for this master
                        if (|master_gnt_vector_addr[m]) begin
                             // Grant active, do not stall based on arb
                        end else begin
                             // No grant yet (Arbitration pending or just lost), must stall
                             // But only if we really requested?
                             // Logic: If requesting (TRANS) and NO GRANT, stall. 
                             HREADYOUT_o[m] = 1'b0;
                        end
                    end
                end
            end
        end
    endgenerate

endmodule
